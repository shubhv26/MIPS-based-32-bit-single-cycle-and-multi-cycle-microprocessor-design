module SQM_CA2_ONES(input logic [3:0]B, 
	            input logic [7:0]A,
	    	    input logic op,  
		    output logic [3:0] Z, 
       		    output logic [7:0]C,
       		    output logic [7:0]Y);
always_comb
begin
reg [7:0]P,Q;
if(op==1'b1)begin
assign C=B*B;
assign Q=C%A;
Y=Q; 
end

else if(op==1'b0)
 begin
P[0]=A[1]?(A[0]?B[3]:B[2]):(A[0]?B[1]:B[0]);
P[1]=A[2]?(A[1]?B[3]:B[2]):(A[1]?B[1]:B[0]);
P[2]=A[3]?(A[2]?B[3]:B[2]):(A[2]?B[1]:B[0]);
P[3]=A[4]?(A[3]?B[3]:B[2]):(A[3]?B[1]:B[0]);
P[4]=A[5]?(A[4]?B[3]:B[2]):(A[4]?B[1]:B[0]);
P[5]=A[6]?(A[5]?B[3]:B[2]):(A[5]?B[1]:B[0]);
P[6]=A[7]?(A[6]?B[3]:B[2]):(A[6]?B[1]:B[0]);
P[7]=A[0]?(A[7]?B[3]:B[2]):(A[7]?B[1]:B[0]);
Y=P;
end

casez(Y)
	8'b11111111 : Z=4'b1000; //8

	8'b11111110 : Z=4'b0111; //7	
	8'b01111111 : Z=4'b0111;

	8'b1111110? : Z=4'b0110; //6
	8'b?0111111 : Z=4'b0110;
	8'b01111110 : Z=4'b0110;
	
	8'b111110?? : Z=4'b0101; //5
	8'b??011111 : Z=4'b0101;
	8'b0111110? : Z=4'b0101;
	8'b?0111110 : Z=4'b0101;

	8'b11110??? : Z=4'b0100; //4
	8'b???01111 : Z=4'b0100;
	8'b011110?? : Z=4'b0100;
	8'b??011110 : Z=4'b0100;
	8'b?011110? : Z=4'b0100;

	8'b1110???0 : Z=4'b0011; //3
	8'b01110??? : Z=4'b0011;
	8'b?01110?? : Z=4'b0011;
	8'b??01110? : Z=4'b0011;
	8'b???01110 : Z=4'b0011;
	8'b0???0111 : Z=4'b0011;
        8'b11100??? : Z=4'b0011;

	8'b110??0?? : Z=4'b0010; //2
	8'b0110??0? : Z=4'b0010;
	8'b?0110??0 : Z=4'b0010;
	8'b??0110?? : Z=4'b0010;
	8'b0??0110? : Z=4'b0010;
	8'b?0??0110 : Z=4'b0010;
	8'b??0??011 : Z=4'b0010;
        8'b?01100?? : Z=4'b0010;

	8'b10?0?0?0 : Z=4'b0001; //1 
	8'b010?0?0? : Z=4'b0001; 
	8'b?010?0?0 : Z=4'b0001; 
	8'b0?010?0? : Z=4'b0001; 
	8'b?0?010?0 : Z=4'b0001; 
	8'b0?0?010? : Z=4'b0001; 
	8'b?0?0?010 : Z=4'b0001; 
	8'b0?0?0?01 : Z=4'b0001;
 
	8'b00000000 : Z=4'b0000; //0
endcase
end
endmodule

